#test1.vhd code
#2024.10.15

