#test2.vhdl code
#2024.10.15

